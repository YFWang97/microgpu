module vga_controller(
    input reset,
    input clk_20,
    input clk_25,
    input vga_data_valid_in,
    input [5:0] vga_data_in,
    output reg vga_ready_out,
    output vsync,
    output hsync,
    output reg [5:0] rgb
);
// Due to the limiation of BRAM on FPGA, only display the central 50 x 50 area
// X index from 180 to 459
// Y index from 100 to 379

localparam X_WINDOW_LOW = 'd295;
localparam X_WINDOW_HIGH = 'd344;
localparam Y_WINDOW_LOW = 'd215;
localparam Y_WINDOW_HIGH = 'd264;

localparam SCREEN_X = 'd799;
localparam SCREEN_Y = 'd524;

reg [5:0] rgb_buf [1:0][2499:0];

reg pingpong;

wire write_buffer;
wire read_buffer;

assign write_buffer = pingpong;
assign read_buffer = ~pingpong; 

reg [9:0] write_x;
reg [9:0] write_y;
reg [11:0] write_index;

wire [9:0] read_x;
wire [9:0] read_y;
reg [11:0] read_index;

wire blank;

always @(posedge clk_25) begin
    if (reset) begin
        pingpong <= 0;
    end
    else begin
        if (vga_ready_out) begin
            pingpong <= ~pingpong;
        end
    end
end

always @(posedge clk_20) begin
    if (vga_data_valid_in) begin
        if ((write_x >= X_WINDOW_LOW && write_x <= X_WINDOW_HIGH) &&
            (write_y >= Y_WINDOW_LOW && write_y <= Y_WINDOW_HIGH)) begin
            rgb_buf[write_buffer][write_index] <= vga_data_in;
        end
    end
end

always @(posedge clk_20) begin
    if (reset) begin
        write_x <= 'd0;
        write_y <= 'd0;
        write_index <= 'd0;
    end
    else begin
        if (vga_data_valid_in) begin
            write_x <= (write_x == 'd799) ? 'd0 : (write_x + 'd1);
            write_y <= (write_x == SCREEN_X) ? ((write_y == SCREEN_Y) ? 'd0 : (write_y + 'd1)) : write_y;
    
            if ((write_x >= X_WINDOW_LOW && write_x <= X_WINDOW_HIGH) &&
                (write_y >= Y_WINDOW_LOW && write_y <= Y_WINDOW_HIGH)) begin
                write_index <= write_index + 'd1;
            end
        end
        else begin
            write_index <= 'd0;
        end
    end
end    

vga v(.clk(clk_25),.reset(reset), .HS (hsync),.VS (vsync), .x (read_x), .y (read_y), .blank (blank));

always @(posedge clk_20) begin
    if (reset) begin
        vga_ready_out <= 0;
    end
    else begin
        if (vga_ready_out) begin
            vga_ready_out <= 0;
        end
        else if (read_x == SCREEN_X && read_y == SCREEN_Y) begin
            vga_ready_out <= 1;
        end
    end
end

always @(posedge clk_25) begin
    if (reset || vga_ready_out) begin
        read_index <= 'd0;
    end
    else begin
        if ((read_x >= X_WINDOW_LOW && read_x <= X_WINDOW_HIGH) &&
            (read_y >= Y_WINDOW_LOW && read_y <= Y_WINDOW_HIGH)) begin
            read_index <= read_index + 'd1;
        end
    end
end

always @(*) begin
    if (blank) rgb = 'd0;
    else if ((read_x >= X_WINDOW_LOW && read_x <= X_WINDOW_HIGH) &&
        (read_y >= Y_WINDOW_LOW && read_y <= Y_WINDOW_HIGH)) begin
        rgb = rgb_buf[read_buffer][read_index];
        //rgb = 6'b101010;
    end
    else begin
        rgb = 6'b010101;
    end
end

endmodule
