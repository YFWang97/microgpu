module dot_product (






);



endmodule
